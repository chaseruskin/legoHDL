--takes all initial library calls from top-level VHD

package template_pkg is

end package;


package body template_pkg is

end package body;