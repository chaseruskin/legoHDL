
package template_pkg is
end package;


package body template_pkg is
end package body;