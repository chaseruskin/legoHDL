--
--Project:
--Author:
--Date:
--Description:
--
library ieee;
use ieee.std_logic_1164.all;

entity template is
    port(
        --list of ports
    );
end entity;


architecture bhv of template is

begin


end architecture;