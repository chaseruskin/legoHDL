--
--  Project:        %PROJECT%
--  Author:         %AUTHOR%
--  Date:           %DATE%
--  Description:
--

library ieee;
use ieee.std_logic_1164.all;

entity template_tb is
end entity;


architecture bhv of template_tb is

begin


end architecture;